`timescale 1ns/10ps 
module MAR
    #(parameter VAL = 0)(
    input wire clk,
    input wire clr,
    input wire [31:0] dIn,
    input wire Rin,
    output reg [8:0] address
);
    always @(posedge clk or negedge clr)
    begin
        if (clr == 0)
            address <= 0;
        else if (Rin)
            address <= dIn[8:0];
    end

    initial
        address = VAL;
endmodule
